module uart_txC 
#(parameter KBAUD = 14'd10416)
(
    input clk,
    input rst, 
    input [7:0] data, 
    input Tx_start, 
    output Tx_done, 
    output Tx_EN, 
    output OUT
);

    
endmodule