module slaveA (
    input ACLK,
    input ARESETn,
    output ARREADY, //read address ready(součástí hand-shaku )
);
    
endmodule