module UartCoder (
    input i_clk,
    input i_reset,
    input i_stb,
    output o_dw_busy,
    input [33:0] i_word,
    output [7:0] out_char
);
    
endmodule