
`ifndef WBDEFS_H

`define WBDEFS_H

`define OPT_UART_RE

`define OPT_SIM = 1

`endif 	//WBDEFS_H