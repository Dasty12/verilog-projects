
`ifndef WBDEFS_H

`define WBDEFS_H

`define OPT_UART_RE



`endif 	//WBDEFS_H