module SPI_top
{
	input clk,
	
};