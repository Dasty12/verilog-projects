module top_osc (
    input clk
);
    




endmodule